-module fpga_cm33
-module led_wf
-module PLL_FREQ
-topmoduleNum 1
-topmodule fpga_cm33
